//============================================================================
//
//  SD card ROM loader and ROM selector for MISTer.
//  Copyright (C) 2019 Kitrinx (aka Rysha)
//
//  Permission is hereby granted, free of charge, to any person obtaining a
//  copy of this software and associated documentation files (the "Software"),
//  to deal in the Software without restriction, including without limitation
//	 the rights to use, copy, modify, merge, publish, distribute, sublicense,
//	 and/or sell copies of the Software, and to permit persons to whom the
//	 Software is furnished to do so, subject to the following conditions:
//
//  The above copyright notice and this permission notice shall be included in
//	 all copies or substantial portions of the Software.
//
//  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
//	 IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
//	 FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
//	 AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
//	 LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
//	 FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
//	 DEALINGS IN THE SOFTWARE.
//
//============================================================================

// Rom layout for Exerion:
// 0x00000 - 0x01FFF = eprom_1 - Background Graphics IC 4B
// 0x02000 - 0x03FFF = eprom_2 - Background Graphics IC 4D
// 0x04000 - 0x05FFF = eprom_3 - Background Graphics IC 4E
// 0x06000 - 0x07FFF = eprom_4 - Background Graphics IC 4H
// 0x08000 - 0x09FFF = eprom_5 - exerion.10 & exerion.11 - Sprites
// 0x0A000 - 0x0BFFF = eprom_6 - exerion.05 - Background Layer Program
// 0x0C000 - 0x0DFFF = eprom_7 - exerion.06 - Foreground Characters
// 0x10000 - 0x15FFF = eprom_8 - eb5 & eb6  - Main Program ROM 1 & 2

module selector
    (
        input logic [24:0] ioctl_addr,
        output logic ep1_cs, ep2_cs, ep3_cs, ep4_cs, ep5_cs, ep6_cs, ep7_cs, ep8_cs
    );

    always_comb begin
        {ep1_cs, ep2_cs, ep3_cs, ep4_cs, ep5_cs, ep6_cs, ep7_cs, ep8_cs} = 0;
        if     (ioctl_addr < 'h2000 ) ep1_cs = 1; // 0x2000 13 - BGL1
        else if(ioctl_addr < 'h04000) ep2_cs = 1; // 0x2000 13 - BGL2
        else if(ioctl_addr < 'h06000) ep3_cs = 1; // 0x2000 13 - BGL3
        else if(ioctl_addr < 'h08000) ep4_cs = 1; // 0x2000 13 - BGL4
        else if(ioctl_addr < 'h0C000) ep5_cs = 1; // 0x4000 14 - Sprites
        else if(ioctl_addr < 'h0e000) ep6_cs = 1; // 0x2000 13 - Background Program
        else if(ioctl_addr < 'h10000) ep7_cs = 1; // 0x2000 13 - Foreground Characters
        else                          ep8_cs = 1; // 0x6000 15 - Main Program //(ioctl_addr < 'h16000)
    end
endmodule

////////////
// EPROMS //
////////////
module eprom_1
    (
        input  logic        CLK,
        input  logic        CLK_DL,
        input  logic        CEN,
        input  logic [12:0] ADDR,
        input  logic [24:0] ADDR_DL,
        input  logic [7:0]  DATA_IN,
        input  logic        CS_DL,
        input  logic        WR,
        output logic [7:0]  DATA
    );

    reg [7:0] DATA_out;
    always @(posedge CLK) DATA <= (CEN) ? 0 : DATA_out;

    dpram_dc #(.widthad_a(13)) eprom_1
             (
                 .clock_a(CLK),
                 .address_a(ADDR[12:0]),
                 .q_a(DATA_out),
                 .clock_b(CLK_DL),
                 .address_b(ADDR_DL[12:0]),
                 .data_b(DATA_IN),
                 .wren_b(WR & CS_DL)
             );
endmodule

module eprom_2
    (
        input  logic        CLK,
        input  logic        CLK_DL,
        input  logic        CEN,
        input  logic [12:0] ADDR,
        input  logic [24:0] ADDR_DL,
        input  logic  [7:0] DATA_IN,
        input  logic        CS_DL,
        input  logic        WR,
        output logic  [7:0] DATA
    );
    reg [7:0] DATA_out;
    always @(posedge CLK) DATA <= (CEN) ? 0 : DATA_out;

    dpram_dc #(.widthad_a(13)) eprom_2
             (
                 .clock_a(CLK),
                 .address_a(ADDR[12:0]),
                 .q_a(DATA_out),
                 .clock_b(CLK_DL),
                 .address_b(ADDR_DL[12:0]),
                 .data_b(DATA_IN),
                 .wren_b(WR & CS_DL)
             );
endmodule

module eprom_3
    (
        input  logic        CLK,
        input  logic        CLK_DL,
        input  logic        CEN,
        input  logic [12:0] ADDR,
        input  logic [24:0] ADDR_DL,
        input  logic  [7:0] DATA_IN,
        input  logic        CS_DL,
        input  logic        WR,
        output logic  [7:0] DATA
    );

    reg [7:0] DATA_out;
    always @(posedge CLK) DATA <= (CEN) ? 0 : DATA_out;

    dpram_dc #(.widthad_a(13)) eprom_3
             (
                 .clock_a(CLK),
                 .address_a(ADDR[12:0]),
                 .q_a(DATA_out),
                 .clock_b(CLK_DL),
                 .address_b(ADDR_DL[12:0]),
                 .data_b(DATA_IN),
                 .wren_b(WR & CS_DL)
             );
endmodule

module eprom_4
    (
        input  logic        CLK,
        input  logic        CLK_DL,
        input  logic        CEN,
        input  logic [12:0] ADDR,
        input  logic [24:0] ADDR_DL,
        input  logic  [7:0] DATA_IN,
        input  logic        CS_DL,
        input  logic        WR,
        output logic  [7:0] DATA
    );
    reg [7:0] DATA_out;
    always @(posedge CLK) DATA <= (CEN) ? 0 : DATA_out;

    dpram_dc #(.widthad_a(13)) eprom_4
             (
                 .clock_a(CLK),
                 .address_a(ADDR[12:0]),
                 .q_a(DATA_out),
                 .clock_b(CLK_DL),
                 .address_b(ADDR_DL[12:0]),
                 .data_b(DATA_IN),
                 .wren_b(WR & CS_DL)
             );
endmodule

module eprom_5
    (
        input  logic        CLK,
        input  logic        CLK_DL,
        input  logic [13:0] ADDR,
        input  logic [24:0] ADDR_DL,
        input  logic  [7:0] DATA_IN,
        input  logic        CS_DL,
        input  logic        WR,
        output logic  [7:0] DATA
    );

    dpram_dc #(.widthad_a(14)) eprom_5
             (
                 .clock_a(CLK),
                 .address_a(ADDR[13:0]),
                 .q_a(DATA[7:0]),

                 .clock_b(CLK_DL),
                 .address_b(ADDR_DL[13:0]),
                 .data_b(DATA_IN),
                 .wren_b(WR & CS_DL)
             );
endmodule

module eprom_6
    (
        input  logic        CLK,
        input  logic        CLK_DL,
        input  logic [12:0] ADDR,
        input  logic [24:0] ADDR_DL,
        input  logic  [7:0] DATA_IN,
        input  logic        CS_DL,
        input  logic        WR,
        output logic  [7:0] DATA
    );

    dpram_dc #(.widthad_a(13)) eprom_6
             (
                 .clock_a(CLK),
                 .address_a(ADDR[12:0]),
                 .q_a(DATA[7:0]),

                 .clock_b(CLK_DL),
                 .address_b(ADDR_DL[12:0]),
                 .data_b(DATA_IN),
                 .wren_b(WR & CS_DL)
             );
endmodule

module eprom_7
    (
        input  logic        CLK,
        input  logic        CLK_DL,
        input  logic [12:0] ADDR,
        input  logic [24:0] ADDR_DL,
        input  logic  [7:0] DATA_IN,
        input  logic        CS_DL,
        input  logic        WR,
        output logic  [7:0] DATA
    );

    dpram_dc #(.widthad_a(13)) eprom_7
             (
                 .clock_a(CLK),
                 .address_a(ADDR[12:0]),
                 .q_a(DATA[7:0]),

                 .clock_b(CLK_DL),
                 .address_b(ADDR_DL[12:0]),
                 .data_b(DATA_IN),
                 .wren_b(WR & CS_DL)
             );
endmodule

module eprom_8
    (
        input  logic        CLK,
        input  logic        CLK_DL,
        input  logic [14:0] ADDR,
        input  logic [24:0] ADDR_DL,
        input  logic  [7:0] DATA_IN,
        input  logic        CS_DL,
        input  logic        WR,
        output logic  [7:0] DATA
    );

    dpram_dc #(.widthad_a(15)) eprom_8
             (
                 .clock_a(CLK),
                 .address_a(ADDR[14:0]),
                 .q_a(DATA[7:0]),

                 .clock_b(CLK_DL),
                 .address_b(ADDR_DL[14:0]),
                 .data_b(DATA_IN),
                 .wren_b(WR & CS_DL)
             );
endmodule

///////////
// PROMS //
///////////
module color_prom_1
    (
        input  logic        CLK,
        input  logic        CLK_DL,
        input  logic  [8:0] ADDR,
        input  logic [24:0] ADDR_DL,
        input  logic  [7:0] DATA_IN,
        input  logic        CS_DL,
        input  logic        WR,
        output logic [ 3:0] DATA
    );

    dpram_dc #(.widthad_a(9)) cprom_1
             (
                 .clock_a(CLK),
                 .address_a(ADDR),
                 .q_a(DATA[3:0]),

                 .clock_b(CLK_DL),
                 .address_b(ADDR_DL[8:0]),
                 .data_b(DATA_IN),
                 .wren_b(WR & CS_DL)
             );
endmodule

module color_prom_2
    (
        input  logic        CLK,
        input  logic        CLK_DL,
        input  logic  [8:0] ADDR,
        input  logic [24:0] ADDR_DL,
        input  logic  [7:0] DATA_IN,
        input  logic        CS_DL,
        input  logic        WR,
        output logic  [3:0] DATA
    );

    dpram_dc #(.widthad_a(9)) cprom_2
             (
                 .clock_a(CLK),
                 .address_a(ADDR),
                 .q_a(DATA[3:0]),

                 .clock_b(CLK_DL),
                 .address_b(ADDR_DL[8:0]),
                 .data_b(DATA_IN),
                 .wren_b(WR & CS_DL)
             );
endmodule

module color_prom_3
    (
        input  logic        CLK,
        input  logic        CLK_DL,
        input  logic  [8:0] ADDR,
        input  logic [24:0] ADDR_DL,
        input  logic  [7:0] DATA_IN,
        input  logic        CS_DL,
        input  logic        WR,
        output logic  [3:0] DATA
    );

    dpram_dc #(.widthad_a(9)) cprom_3
             (
                 .clock_a(CLK),
                 .address_a(ADDR),
                 .q_a(DATA[3:0]),

                 .clock_b(CLK_DL),
                 .address_b(ADDR_DL[8:0]),
                 .data_b(DATA_IN),
                 .wren_b(WR & CS_DL)
             );
endmodule
